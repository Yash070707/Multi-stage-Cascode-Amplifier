magic
tech scmos
timestamp 1668071664
<< nwell >>
rect -42 -457 95 184
<< ntransistor >>
rect 2 -524 6 -492
rect 2 -581 6 -555
<< ptransistor >>
rect 2 -81 6 135
rect 2 -426 6 -128
<< ndiffusion >>
rect -5 -493 2 -492
rect -1 -497 2 -493
rect -5 -524 2 -497
rect 6 -493 13 -492
rect 6 -497 9 -493
rect 6 -524 13 -497
rect -5 -558 2 -555
rect -1 -562 2 -558
rect -5 -581 2 -562
rect 6 -558 13 -555
rect 6 -562 9 -558
rect 6 -581 13 -562
<< pdiffusion >>
rect -5 125 2 135
rect -1 121 2 125
rect -5 -81 2 121
rect 6 89 13 135
rect 6 85 9 89
rect 6 -81 13 85
rect -5 -149 2 -128
rect -1 -153 2 -149
rect -5 -426 2 -153
rect 6 -149 13 -128
rect 6 -153 9 -149
rect 6 -426 13 -153
<< ndcontact >>
rect -5 -497 -1 -493
rect 9 -497 13 -493
rect -5 -562 -1 -558
rect 9 -562 13 -558
<< pdcontact >>
rect -5 121 -1 125
rect 9 85 13 89
rect -5 -153 -1 -149
rect 9 -153 13 -149
<< psubstratepcontact >>
rect -22 -603 -18 -599
rect 0 -603 4 -599
rect 25 -603 29 -599
<< nsubstratencontact >>
rect -25 157 -21 161
rect 1 157 5 161
rect 22 157 26 161
<< polysilicon >>
rect 2 137 4 142
rect 2 135 6 137
rect 2 -85 6 -81
rect 4 -126 6 -121
rect 2 -128 6 -126
rect 2 -430 6 -426
rect 2 -490 4 -485
rect 2 -492 6 -490
rect 2 -528 6 -524
rect 2 -553 4 -548
rect 2 -555 6 -553
rect 2 -585 6 -581
<< polycontact >>
rect 4 137 8 142
rect 0 -126 4 -121
rect 4 -490 8 -485
rect 4 -553 8 -548
<< metal1 >>
rect -33 161 42 164
rect -33 157 -25 161
rect -21 157 1 161
rect 5 157 22 161
rect 26 157 42 161
rect -33 154 42 157
rect -25 125 -21 154
rect 8 137 12 142
rect -25 121 -5 125
rect 13 85 38 89
rect -4 -126 0 -121
rect 34 -149 38 85
rect -25 -153 -5 -149
rect 13 -153 38 -149
rect -25 -465 -21 -153
rect -25 -469 -4 -465
rect -25 -493 -21 -469
rect 8 -490 13 -485
rect -25 -497 -5 -493
rect 13 -497 30 -493
rect 8 -553 13 -548
rect 26 -558 30 -497
rect -22 -562 -5 -558
rect 13 -562 30 -558
rect -22 -594 -18 -562
rect -31 -599 47 -594
rect -31 -603 -22 -599
rect -18 -603 0 -599
rect 4 -603 25 -599
rect 29 -603 47 -599
rect -31 -608 47 -603
<< labels >>
rlabel metal1 -1 159 -1 159 1 vdd!
rlabel metal1 -11 -601 -11 -601 1 gnd!
rlabel metal1 -2 -124 -2 -124 1 Vbias2
rlabel metal1 10 140 10 140 1 Vbias1
rlabel metal1 10 -487 10 -487 1 Vbias3
rlabel metal1 10 -550 10 -550 1 Vinput
rlabel metal1 36 -42 36 -42 1 w1
rlabel metal1 28 -524 28 -524 1 w3
rlabel metal1 -8 -467 -8 -467 1 Vout
<< end >>
